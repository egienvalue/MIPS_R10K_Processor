//*****************************************************************************
// Filename: core.v
// Discription: core top level integration, instantiate new feature modules
// 				here
// Author: group 5
// Version History
//   <11/5> initial creation: integrate without br_stack, br_predictor, LSQ
//*****************************************************************************
`timescale 1ns/100ps

module core (
		input									clk,
		input									rst,

		input			[3:0]					mem2proc_response,
		input			[63:0]					mem2proc_data,
		input			[3:0]					mem2proc_tag,
	
		output	logic	[1:0]					proc2mem_command,
		output	logic	[63:0]					proc2mem_addr,
		output	logic	[63:0]					proc2mem_data,




	);



	//---------------------------------------------------------------
	// signals for Icache
	//---------------------------------------------------------------


	//---------------------------------------------------------------
	// signals for if_stage
	//---------------------------------------------------------------
	
	
	//---------------------------------------------------------------
	// signals for branch predictor
	//---------------------------------------------------------------


	//---------------------------------------------------------------
	// signals for dispatch
	//---------------------------------------------------------------


	//---------------------------------------------------------------
	// signals for rs
	//---------------------------------------------------------------


	//---------------------------------------------------------------
	// signals for rob
	//---------------------------------------------------------------


	//---------------------------------------------------------------
	// signals for map table and free list
	//---------------------------------------------------------------


	//---------------------------------------------------------------
	// signals for fu
	//---------------------------------------------------------------


	//---------------------------------------------------------------
	// signals for early branch recovery (br stack)
	//---------------------------------------------------------------
	

	//---------------------------------------------------------------
	// signals for LSQ
	//---------------------------------------------------------------
	
	
	//---------------------------------------------------------------
	// signals for Dcache
	//---------------------------------------------------------------
	
	

	//===============================================================
	// Icache instantiation
	//===============================================================
	

	//===============================================================
	// if_stage instantiation
	//===============================================================
	if_stage(
				  .clk,                      // system clk
				  .rst,                      // system rst
				  					        // makes pipeline behave as single-cycle
				  .branch_i,
				  .br_dirp_i,
				  .return_i,
				  .ras_target_i,
				  .br_predict_target_PC_i,
				  .br_flush_target_PC_i,
				  .Imem2proc_data,		        // Data coming back from instruction-memory
				  .Imem_valid,
				  .br_flush_en_i,
				  .id_request_i,

				  .proc2Imem_addr,		// Address sent to Instruction memory
				  .if_NPC_out,			// PC of instruction after fetched (PC+4).
				  .if_IR_out,			// fetched instruction out
				  .if_valid_inst_out	    // when low, instruction is garbage
				  //output logic		  if2id_empty_o
           );


	//===============================================================
	// branch predictor instantiation
	//===============================================================
	

	//===============================================================
	// dispatch instantiation
	//===============================================================
	

	//===============================================================
	// rs instantiation
	//===============================================================
	

	//===============================================================
	// map table and free list instantiation
	//===============================================================
	

	//===============================================================
	// fu instantiation
	//===============================================================
		

	//===============================================================
	// early branch recovery instantiation
	//===============================================================
	

	//===============================================================
	// LSQ instantiation
	//===============================================================
	

	//===============================================================
	// Dcache instantiation
	//===============================================================
	


