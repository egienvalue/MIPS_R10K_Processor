
`define SD                         #1
`define CLK_PERIOD                 #1000
`define CLK_PERIOD_HALF            #500

