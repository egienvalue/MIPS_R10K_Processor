// ****************************************************************************
// Filename: alu2.v
// Discription: alu for branch condition calculation
// Author: Jun
// Version History:
// 	intial creation: 10/26/2017
// 	***************************************************************************
module alu1 (

		input		[63:0] br_disp_i;
		input		[63:0] npc;
		input				
		
	
		);
